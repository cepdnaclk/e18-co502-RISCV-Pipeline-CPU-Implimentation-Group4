// Advanced Computer Architecture (CO502)
// Design: ID_EX Pipeline Register
// Group Number: 4
// E Numbers: E/18/077, E/18/397, E/18/402
// Names: Nipun Dharmarathne, Shamod Wijerathne, Chatura Wimalasiri 

module ID_EX_register(
	CLK,
	RESET,
	WRITE_ENABLE_IN,
	MUXDATAMEM_SELECT_IN,
	MEM_READ_IN,
	MEM_WRITE_IN,
	MUXJAL_SELECT_IN,
	ALUOP_IN,
	MUXIMM_SELECT_IN,
	MUXPC_SELECT_IN,
	BRANCH_IN,
	JUMP_IN,
	PC_DIRECT_OUT_IN,
	SIGN_ZERO_EXTEND,
	PC_PLUS_4_OUT_IN,
	OUT1_IN,
	OUT2_IN,
	RD_IN,
	FUNCT3_IN,
	WRITE_ENABLE_OUT,
	MUXDATAMEM_SELECT_OUT,
	MEM_READ_OUT,
	MEM_WRITE_OUT,
	MUXJAL_SELECT_OUT,
	ALUOP_OUT,
	MUXIMM_SELECT_OUT,
	MUXPC_SELECT_OUT,
	BRANCH_OUT,
	JUMP_OUT,
	PC_DIRECT_OUT_OUT,
	SIGN_ZERO_EXTEND_OUT,
	PC_PLUS_4_OUT_OUT,
	OUT1_OUT,
	OUT2_OUT,
	RD_OUT,
	FUNCT3_OUT,
	BUSYWAIT
);
	
	//port declarations
	input CLK, RESET, WRITE_ENABLE_IN, MUXDATAMEM_SELECT_IN, MEM_READ_IN, MEM_WRITE_IN, MUXJAL_SELECT_IN, MUXIMM_SELECT_IN, MUXPC_SELECT_IN, BRANCH_IN, JUMP_IN, BUSYWAIT;
	input [2:0] FUNCT3_IN;
	input [4:0] ALUOP_IN, RD_IN;
	input [31:0] PC_DIRECT_OUT_IN, SIGN_ZERO_EXTEND, PC_PLUS_4_OUT_IN, OUT1_IN, OUT2_IN;
	
	output reg WRITE_ENABLE_OUT, MUXDATAMEM_SELECT_OUT, MEM_READ_OUT, MEM_WRITE_OUT, MUXJAL_SELECT_OUT, MUXIMM_SELECT_OUT, MUXPC_SELECT_OUT, BRANCH_OUT, JUMP_OUT;
	output reg [2:0] FUNCT3_OUT;
	output reg [4:0] ALUOP_OUT, RD_OUT;
	output reg [31:0] PC_DIRECT_OUT_OUT, SIGN_ZERO_EXTEND_OUT, PC_PLUS_4_OUT_OUT, OUT1_OUT, OUT2_OUT;
	
	
	// reset the registers
	always @ (*) begin
        if (RESET) begin
			#1
			WRITE_ENABLE_OUT = 1'dx; 
			MUXDATAMEM_SELECT_OUT = 1'dx; 
			MEM_READ_OUT = 1'dx; 
			MEM_WRITE_OUT = 1'dx; 
			MUXJAL_SELECT_OUT = 1'dx; 
			MUXIMM_SELECT_OUT = 1'dx; 
			MUXPC_SELECT_OUT = 1'dx; 
			BRANCH_OUT = 1'dx; 
			JUMP_OUT = 1'dx; 
			
			FUNCT3_OUT = 3'dx;
			
			ALUOP_OUT = 5'dx;
			RD_OUT = 5'dx;
			
			PC_DIRECT_OUT_OUT = 32'dx;
			SIGN_ZERO_EXTEND_OUT = 32'dx;
			PC_PLUS_4_OUT_OUT = 32'dx;
			OUT1_OUT = 32'dx;
			OUT2_OUT = 32'dx;
		end
	end
	
	
	// input data tranmits to outputs at the positive edge of the clock
	// At this moment, reset must be low
	// Assignments to outputs happen simultaneously
	always @ (posedge CLK) begin
        if (!BUSYWAIT && !RESET) begin
			#1
			WRITE_ENABLE_OUT <= WRITE_ENABLE_IN;
			MUXDATAMEM_SELECT_OUT <= MUXDATAMEM_SELECT_IN;
			MEM_READ_OUT <= MEM_READ_IN;
			MEM_WRITE_OUT <= MEM_WRITE_IN;
			MUXJAL_SELECT_OUT <= MUXJAL_SELECT_IN;
			MUXIMM_SELECT_OUT <= MUXIMM_SELECT_IN;
			MUXPC_SELECT_OUT <= MUXPC_SELECT_IN;
			BRANCH_OUT <= BRANCH_IN;
			JUMP_OUT <= JUMP_IN;
			
			FUNCT3_OUT <= FUNCT3_IN;
			
			ALUOP_OUT <= ALUOP_IN;
			RD_OUT <= RD_IN;
			
			PC_DIRECT_OUT_OUT <= PC_DIRECT_OUT_IN;
			SIGN_ZERO_EXTEND_OUT <= SIGN_ZERO_EXTEND;
			PC_PLUS_4_OUT_OUT <= PC_PLUS_4_OUT_IN;
			OUT1_OUT <= OUT1_IN;
			OUT2_OUT <= OUT2_IN;
		
		
		end
	end

endmodule
	
	
	
	
	