`timescale  1ns/100ps

`include "../RegisterFile/reg_file.v"
`include "../Sign_Zero_Extend/Sign_Zero_Extend.v"
`include "../ControlUnit/control_unit.v"

`include "../Pipeline_Registers/2_ID_EX/ID_EX_register.v"

`include "../Other_modules/mux_2x1_32bit/mux_2x1_32bit.v"
`include "../ALU/alu.v"
`include "../Jump_Controller/Jump_Controller.v"
`include "../Pipeline_Registers/3_EX_MEM/EX_MEM_register.v"

`include "../Data_Memory/Data_Cache.v"
`include "../Data_Memory/Data_Memory.v"
`include "../Pipeline_Registers/4_MEM_WB/MEM_WB_register.v"

`include "../Adder_32bit_plus4/adder_32bit_plus_4.v"
`include "pc.v"
`include "../InstructionMemory/instruction_cache.v"
`include "../InstructionMemory/instruction_memory.v"
`include "../Pipeline_Registers/1_IF_ID/IF_ID_register.v"

module cpu(CLK, RESET);
// port declaration
input RESET, CLK; 

wire WRITE_REG, MUXPC_SELECT, MUXIMM_SELECT, MUXJAL_SELECT, MUXDATAMEM_SELECT, WRITE_ENABLE, MEM_READ, MEM_WRITE, BRANCH, JUMP;
wire [31:0] INSTRUCTION, IN_REG, OUT1_REG, OUT2_REG, SIGN_ZERO_EXTEND,  PC_DIRECT_OUT_IN, PC_PLUS_4_OUT_IN;
wire [4:0] MEM_WB_INADDRESS, ALUOP;
wire[2:0] MUXIMMTYPE_SELECT;

// ID/EX and EX/MEM stage wires
wire EQ_FLAG, LT_FLAG, LTU_FLAG, PC_MUX_CONTROL, REG_FLUSH;
wire [31:0] DATA1, DATA2, RESULT_ALU, MUXJAL_OUT, BRANCH_OR_JUMP_ADDR;

// EX/MEM and MEM/WB stage wires
wire MEM_BUSYWAIT, MEM_MEM_READ, MEM_MEM_WRITE; 
wire [27:0] MEM_BLOCK_ADDR;
wire [31:0] CACHE_READ_OUT;
wire [127:0] DATA_MEM_READ_OUT, DATA_MEM_WRITE_OUT;

// MEM/WB and IF/ID stage
wire [31:0] PC, PC_PLUS_4, PC_MUX_OUT;


// ID_EX Register Outputs
wire WRITE_ENABLE_OUT, MUXDATAMEM_SELECT_OUT, MEM_READ_OUT, MEM_WRITE_OUT, MUXJAL_SELECT_OUT, MUXIMM_SELECT_OUT, MUXPC_SELECT_OUT, BRANCH_OUT, JUMP_OUT;
wire [2:0] FUNCT3_OUT;
wire [4:0] ALUOP_OUT, RD_OUT;
wire [31:0] PC_DIRECT_OUT_OUT, SIGN_ZERO_EXTEND_OUT, PC_PLUS_4_OUT_OUT, OUT1_OUT, OUT2_OUT;

// EX_MEM Register Outputs
wire WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, MEM_READ_OUT_EX_MEM, MEM_WRITE_OUT_EX_MEM;
wire [2:0] FUNCT3_OUT_EX_MEM;
wire [4:0] RD_OUT_EX_MEM;
wire [31:0] MUXJAL_OUT_EX_MEM, OUT2_OUT_EX_MEM;

// MEM_WB Register Outputs
wire  MUXDATAMEM_SELECT_OUT_MEM_WB;
wire [31:0] CACHE_READ_OUT_MEM_WB, MUXJAL_OUT_MEM_WB;

wire [31:0] READINST;
wire [27:0] MEM_ADDRESS_TO_CACHE;
wire [127:0] MEM_READINST;
wire I_BUSYWAIT, I_MEM_READ, I_MEM_BUSYWAIT;

wire BUSYWAIT, D_BUSYWAIT;

assign BUSYWAIT = D_BUSYWAIT || I_BUSYWAIT;

/* 
	IF/ID and ID/EX stage
*/
reg_file myreg(IN_REG, OUT1_REG, OUT2_REG, MEM_WB_INADDRESS, INSTRUCTION[19:15], INSTRUCTION[24:20], WRITE_REG, CLK, RESET); 
control_unit mycu(INSTRUCTION, ALUOP,  MUXIMMTYPE_SELECT, MUXPC_SELECT, MUXIMM_SELECT, MUXJAL_SELECT, MUXDATAMEM_SELECT, WRITE_ENABLE, MEM_READ, MEM_WRITE, BRANCH, JUMP);
Sign_Zero_Extend signZeroExtend(INSTRUCTION,MUXIMMTYPE_SELECT, SIGN_ZERO_EXTEND );
ID_EX_register myIDEX(CLK,REG_FLUSH,WRITE_ENABLE,MUXDATAMEM_SELECT,MEM_READ,MEM_WRITE,MUXJAL_SELECT,ALUOP,MUXIMM_SELECT,MUXPC_SELECT,BRANCH,JUMP,PC_DIRECT_OUT_IN,SIGN_ZERO_EXTEND,PC_PLUS_4_OUT_IN,OUT1_REG,OUT2_REG, INSTRUCTION[11:7],INSTRUCTION[14:12],
WRITE_ENABLE_OUT,MUXDATAMEM_SELECT_OUT,MEM_READ_OUT,MEM_WRITE_OUT,MUXJAL_SELECT_OUT,ALUOP_OUT,MUXIMM_SELECT_OUT,MUXPC_SELECT_OUT,BRANCH_OUT,JUMP_OUT,PC_DIRECT_OUT_OUT,SIGN_ZERO_EXTEND_OUT,PC_PLUS_4_OUT_OUT,OUT1_OUT,OUT2_OUT,RD_OUT,FUNCT3_OUT,BUSYWAIT);

/* 
	ID/EX and EX/MEM stage
*/
mux_2x1_32bit muxpc(OUT1_OUT, PC_DIRECT_OUT_OUT, DATA1, MUXPC_SELECT_OUT);
mux_2x1_32bit muximm(OUT2_OUT, SIGN_ZERO_EXTEND_OUT, DATA2, MUXIMM_SELECT_OUT);
alu myalu(DATA1, DATA2, RESULT_ALU, ALUOP_OUT, EQ_FLAG, LT_FLAG, LTU_FLAG);
mux_2x1_32bit muxjal(RESULT_ALU, PC_PLUS_4_OUT_OUT, MUXJAL_OUT, MUXJAL_SELECT_OUT);
Jump_Controller myjump_controller(RESULT_ALU, SIGN_ZERO_EXTEND_OUT, FUNCT3_OUT, BRANCH_OUT, JUMP_OUT, EQ_FLAG, LT_FLAG, LTU_FLAG, BRANCH_OR_JUMP_ADDR, PC_MUX_CONTROL, REG_FLUSH);

EX_MEM_register my_ex_mem_register(CLK, REG_FLUSH, WRITE_ENABLE_OUT, MUXDATAMEM_SELECT_OUT, MEM_READ_OUT, MEM_WRITE_OUT, MUXJAL_OUT, OUT2_OUT, RD_OUT, FUNCT3_OUT, 
 WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, MEM_READ_OUT_EX_MEM, MEM_WRITE_OUT_EX_MEM, MUXJAL_OUT_EX_MEM, OUT2_OUT_EX_MEM, RD_OUT_EX_MEM, FUNCT3_OUT_EX_MEM, BUSYWAIT);



/* 
	EX/MEM and MEM/WB stage
*/
dcache my_data_cache(CLK, RESET, MEM_READ_OUT_EX_MEM, MEM_WRITE_OUT_EX_MEM, MUXJAL_OUT_EX_MEM, OUT2_OUT_EX_MEM, MEM_BUSYWAIT, DATA_MEM_READ_OUT, CACHE_READ_OUT, MEM_MEM_READ, MEM_MEM_WRITE, D_BUSYWAIT, MEM_BLOCK_ADDR, DATA_MEM_WRITE_OUT);
data_memory my_data_memory(CLK, RESET, MEM_MEM_READ, MEM_MEM_WRITE, MEM_BLOCK_ADDR, DATA_MEM_WRITE_OUT, DATA_MEM_READ_OUT, MEM_BUSYWAIT);

MEM_WB_register my_mem_wb_register(CLK, REG_FLUSH, WRITE_ENABLE_OUT_EX_MEM,  MUXDATAMEM_SELECT_OUT_EX_MEM, CACHE_READ_OUT, MUXJAL_OUT_EX_MEM, RD_OUT_EX_MEM, 
	WRITE_REG, MUXDATAMEM_SELECT_OUT_MEM_WB, CACHE_READ_OUT_MEM_WB, MUXJAL_OUT_MEM_WB, MEM_WB_INADDRESS, BUSYWAIT);

/* 
	MEM/WB and IF/ID stage
*/
mux_2x1_32bit muxdatamem(MUXJAL_OUT_MEM_WB, CACHE_READ_OUT_MEM_WB, IN_REG, MUXDATAMEM_SELECT_OUT_EX_MEM);


mux_2x1_32bit pc_mux(PC_PLUS_4, BRANCH_OR_JUMP_ADDR, PC_MUX_OUT, PC_MUX_CONTROL);
pc_module my_pc(PC_MUX_OUT, PC, RESET, CLK, BUSYWAIT);
adder_32bit_plus_4 my_adder_32bit_plus_4(PC, PC_PLUS_4);


instruction_cache my_instruction_cache(CLK,RESET, PC, READINST,   I_BUSYWAIT, MEM_ADDRESS_TO_CACHE, I_MEM_READ, MEM_READINST, I_MEM_BUSYWAIT);

instruction_memory my_instruction_memory( CLK,I_MEM_READ,MEM_ADDRESS_TO_CACHE,MEM_READINST,I_MEM_BUSYWAIT);

IF_ID_register myIFID(CLK,REG_FLUSH,READINST,PC_PLUS_4,PC,INSTRUCTION,PC_PLUS_4_OUT_IN,PC_DIRECT_OUT_IN,BUSYWAIT);


endmodule